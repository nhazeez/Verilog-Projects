program testcase();
   import uvm_pkg::*;

   `include "testclass.sv"

   initial begin
      run_test();
   end
endprogram
